`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/24/2023 02:27:45 PM
// Design Name: 
// Module Name: PC
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


// module PC(
//     input clk,
//     input [7:0] PC_in,
//     output[7:0] PC_out
//     );
//     reg [7:0] out;
//     assign PC_out = out;
//     initial out = 8'd0;
//     always@(posedge clk)
//         out <= PC_in;
// endmodule
